
module test(
	input wire a,
	output wire b
);

	parameter sp = 5'd29;
	assign b = sp;
endmodule