module mux_PC_memory (
    input wire selector,
    input wire [31:0] Data_0;
    input wire [31:0] Data_1;
);
    
endmodule